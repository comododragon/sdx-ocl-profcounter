`ifndef COMMANDS_VH
`define COMMANDS_VH

`define COMM_NOP 'h0
`define COMM_STAMP 'h1
`define COMM_HOLD 'h2
`define COMM_FINISH 'h3

`endif
