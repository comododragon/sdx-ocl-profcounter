`ifndef COMMANDS_VH
`define COMMANDS_VH

`define COMM_NOP 'h0
`define COMM_STAMP 'hD
`define COMM_HOLD 'hE
`define COMM_FINISH 'hF

`endif
